module clk(
    input wire clk
);

endmodule