module clock(
    input clk
);

endmodule 