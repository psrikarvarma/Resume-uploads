module clock(input wire clk);

endmodule 